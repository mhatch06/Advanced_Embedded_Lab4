----------------------------------------------------------------------------------

----------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE work.hdmi_package.ALL;
PACKAGE acquireToHDMI_package IS
  -- Clock period definitions
  CONSTANT clk_period : TIME := 20 ns; -- 50Mhz crystal input (XTL_IN).

  -- You need to complete this
  TYPE state_type IS (RESET_STATE);
  ---------------------------- CONTROL WORD -----------------------------
  CONSTANT CW_WIDTH : NATURAL := 22;
  CONSTANT CONTROL_CW_WIDTH : NATURAL := xx;

  CONSTANT CLEAR_STORE_FLAG_CW_BIT_INDEX : NATURAL := 21;
  CONSTANT SET_STORE_FLAG_CW_BIT_INDEX : NATURAL := 20;
  CONSTANT TRIG_CH2_WRITE_CW_BIT_INDEX : NATURAL := 19;
  CONSTANT TRIG_CH1_WRITE_CW_BIT_INDEX : NATURAL := 18;
  CONSTANT CONVERSION_PLUS_READOUT_CW_BIT_INDEX : NATURAL := 17;
  CONSTANT SAMPLE_TIMER_ROLLOVER_CW_BIT_INDEX : NATURAL := 16;
  CONSTANT DATA_STORAGE_CH2_WRITE_CW_BIT_INDEX : NATURAL := 15;
  CONSTANT DATA_STORAGE_CH1_WRITE_CW_BIT_INDEX : NATURAL := 14;
  CONSTANT CONVST_CW_BIT_INDEX : NATURAL := 13;
  CONSTANT RD_CW_BIT_INDEX : NATURAL := 12;
  CONSTANT CS_CW_BIT_INDEX : NATURAL := 11;
  CONSTANT RESET_AD76076_CW_BIT_INDEX : NATURAL := 10;
  CONSTANT DATA_STORAGE_COUNTER_CW_BIT1_INDEX : NATURAL := 9;
  CONSTANT DATA_STORAGE_COUNTER_CW_BIT0_INDEX : NATURAL := 8;
  CONSTANT SAMPLING_COUNTER_CW_BIT1_INDEX : NATURAL := 7;
  CONSTANT SAMPLING_COUNTER_CW_BIT0_INDEX : NATURAL := 6;
  CONSTANT SAMPLING_RATE_SELECT_CW_BIT1_INDEX : NATURAL := 5;
  CONSTANT SAMPLING_RATE_SELECT_CW_BIT0_INDEX : NATURAL := 4;
  CONSTANT LONG_DELAY_COUNTER_CW_BIT1_INDEX : NATURAL := 3;
  CONSTANT LONG_DELAY_COUNTER_CW_BIT0_INDEX : NATURAL := 2;
  CONSTANT SHORT_DELAY_COUNTER_CW_BIT1_INDEX : NATURAL := 1;
  CONSTANT SHORT_DELAY_COUNTER_CW_BIT0_INDEX : NATURAL := 0;

  ---------------------------- STATUS WORD -----------------------------
  CONSTANT SW_WIDTH : NATURAL := 12;
  CONSTANT DATAPATH_SW_WIDTH : NATURAL := 6;

  CONSTANT AD7606_BUSY_SW_INDEX : NATURAL := 11;
  CONSTANT STORE_TO_BRAM_SW_INDEX : NATURAL := 10;
  CONSTANT CH2_TRIGGER_SW_INDEX : NATURAL := 9;
  CONSTANT CH1_TRIGGER_SW_INDEX : NATURAL := 8;
  CONSTANT LONG_DELAY_SW_INDEX : NATURAL := 7;
  CONSTANT SHORT_DELAY_SW_INDEX : NATURAL := 6;
  CONSTANT FULL_SW_INDEX : NATURAL := 5;
  CONSTANT SAMPLE_SW_INDEX : NATURAL := 4;
  CONSTANT TRIGGER_SW_INDEX : NATURAL := 3;
  CONSTANT STORE_SW_INDEX : NATURAL := 2;
  CONSTANT FORCED_SW_INDEX : NATURAL := 1;
  CONSTANT SINGLE_SW_INDEX : NATURAL := 0;
  ------------------------- OTHER CONSTANTS ----------------------------

  CONSTANT LONG_DELAY_50Mhz_CONST_WIDTH : NATURAL := 24;
  CONSTANT LONG_DELAY_50Mhz_COUNTS : STD_LOGIC_VECTOR(LONG_DELAY_50Mhz_CONST_WIDTH - 1 DOWNTO 0) := x"00FFFF";

  CONSTANT SHORT_DELAY_50Mhz_CONST_WIDTH : NATURAL := 8;
  CONSTANT SHORT_DELAY_50Mhz_COUNTS : STD_LOGIC_VECTOR(SHORT_DELAY_50Mhz_CONST_WIDTH - 1 DOWNTO 0) := x"10";

  CONSTANT HIGHEST_RATE : STD_LOGIC_VECTOR(31 DOWNTO 0) := STD_LOGIC_VECTOR(to_unsigned(300, 32));
  CONSTANT HIGH_RATE : STD_LOGIC_VECTOR(31 DOWNTO 0) := STD_LOGIC_VECTOR(to_unsigned(600, 32));
  CONSTANT LOWEST_RATE : STD_LOGIC_VECTOR(31 DOWNTO 0) := STD_LOGIC_VECTOR(to_unsigned(1200, 32));
  CONSTANT LOW_RATE : STD_LOGIC_VECTOR(31 DOWNTO 0) := STD_LOGIC_VECTOR(to_unsigned(2400, 32));
  -----------------------------  HDMI  --------------------------------

  CONSTANT VIDEO_WIDTH_IN_BITS : NATURAL := 11; -- 1650 "pixels" wide, this include FP, SYNCH and BP

  CONSTANT H_ACTIVE : STD_LOGIC_VECTOR(VIDEO_WIDTH_IN_BITS - 1 DOWNTO 0) := STD_LOGIC_VECTOR(to_unsigned(1280, VIDEO_WIDTH_IN_BITS));
  CONSTANT H_FP : STD_LOGIC_VECTOR(VIDEO_WIDTH_IN_BITS - 1 DOWNTO 0) := STD_LOGIC_VECTOR(to_unsigned(110, VIDEO_WIDTH_IN_BITS));
  CONSTANT H_SYNC : STD_LOGIC_VECTOR(VIDEO_WIDTH_IN_BITS - 1 DOWNTO 0) := STD_LOGIC_VECTOR(to_unsigned(40, VIDEO_WIDTH_IN_BITS));
  CONSTANT H_BP : STD_LOGIC_VECTOR(VIDEO_WIDTH_IN_BITS - 1 DOWNTO 0) := STD_LOGIC_VECTOR(to_unsigned(220, VIDEO_WIDTH_IN_BITS));

  CONSTANT H_NOTACTIVE : STD_LOGIC_VECTOR(VIDEO_WIDTH_IN_BITS - 1 DOWNTO 0) := H_FP + H_SYNC + H_BP;
  CONSTANT H_TOTAL : STD_LOGIC_VECTOR(VIDEO_WIDTH_IN_BITS - 1 DOWNTO 0) := H_ACTIVE + H_FP + H_SYNC + H_BP;

  CONSTANT V_ACTIVE : STD_LOGIC_VECTOR(VIDEO_WIDTH_IN_BITS - 1 DOWNTO 0) := STD_LOGIC_VECTOR(to_unsigned(720, VIDEO_WIDTH_IN_BITS));
  CONSTANT V_FP : STD_LOGIC_VECTOR(VIDEO_WIDTH_IN_BITS - 1 DOWNTO 0) := STD_LOGIC_VECTOR(to_unsigned(5, VIDEO_WIDTH_IN_BITS));
  CONSTANT V_SYNC : STD_LOGIC_VECTOR(VIDEO_WIDTH_IN_BITS - 1 DOWNTO 0) := STD_LOGIC_VECTOR(to_unsigned(5, VIDEO_WIDTH_IN_BITS));
  CONSTANT V_BP : STD_LOGIC_VECTOR(VIDEO_WIDTH_IN_BITS - 1 DOWNTO 0) := STD_LOGIC_VECTOR(to_unsigned(20, VIDEO_WIDTH_IN_BITS));

  CONSTANT V_TOTAL : STD_LOGIC_VECTOR(VIDEO_WIDTH_IN_BITS - 1 DOWNTO 0) := V_ACTIVE + V_FP + V_SYNC + V_BP;
  -- You should create constants for your display so that you can easily move the
  -- oscilloscope face around the display.  This makes it easier to make things look
  -- just right
  -- Finish and add more 
  CONSTANT L_EDGE : STD_LOGIC_VECTOR(VIDEO_WIDTH_IN_BITS - 1 DOWNTO 0) := STD_LOGIC_VECTOR(to_unsigned(139, VIDEO_WIDTH_IN_BITS));
  CONSTANT R_EDGE : STD_LOGIC_VECTOR(VIDEO_WIDTH_IN_BITS - 1 DOWNTO 0) := STD_LOGIC_VECTOR(to_unsigned(1139, VIDEO_WIDTH_IN_BITS));
  CONSTANT WIDTH : STD_LOGIC_VECTOR(VIDEO_WIDTH_IN_BITS - 1 DOWNTO 0) := STD_LOGIC_VECTOR(to_unsigned(5, VIDEO_WIDTH_IN_BITS));

  CONSTANT T_EDGE : STD_LOGIC_VECTOR(VIDEO_WIDTH_IN_BITS - 1 DOWNTO 0) := STD_LOGIC_VECTOR(to_unsigned(59, VIDEO_WIDTH_IN_BITS));
  CONSTANT B_EDGE : STD_LOGIC_VECTOR(VIDEO_WIDTH_IN_BITS - 1 DOWNTO 0) := STD_LOGIC_VECTOR(to_unsigned(659, VIDEO_WIDTH_IN_BITS));

  CONSTANT H_HATCH : STD_LOGIC_VECTOR(VIDEO_WIDTH_IN_BITS - 1 DOWNTO 0) := STD_LOGIC_VECTOR(to_unsigned(359, VIDEO_WIDTH_IN_BITS));
  CONSTANT V_HATCH : STD_LOGIC_VECTOR(VIDEO_WIDTH_IN_BITS - 1 DOWNTO 0) := STD_LOGIC_VECTOR(to_unsigned(639, VIDEO_WIDTH_IN_BITS));

  -- You should create constants for your display colors so that modify the colors 
  -- to make things look just right.
  CONSTANT BORDER_R : STD_LOGIC_VECTOR(7 DOWNTO 0) := X"FF";
  CONSTANT BORDER_G : STD_LOGIC_VECTOR(7 DOWNTO 0) := X"FF";
  CONSTANT BORDER_B : STD_LOGIC_VECTOR(7 DOWNTO 0) := X"FF";

  -- Finish and add more 
  CONSTANT GRID_R : STD_LOGIC_VECTOR(7 DOWNTO 0) := X"40";
  CONSTANT GRID_G : STD_LOGIC_VECTOR(7 DOWNTO 0) := X"40";
  CONSTANT GRID_B : STD_LOGIC_VECTOR(7 DOWNTO 0) := X"40";

  CONSTANT TRIG_R : STD_LOGIC_VECTOR(7 DOWNTO 0) := X"00";
  CONSTANT TRIG_G : STD_LOGIC_VECTOR(7 DOWNTO 0) := X"FF";
  CONSTANT TRIG_B : STD_LOGIC_VECTOR(7 DOWNTO 0) := X"FF";

  CONSTANT CH1_R : STD_LOGIC_VECTOR(7 DOWNTO 0) := X"FF";
  CONSTANT CH1_G : STD_LOGIC_VECTOR(7 DOWNTO 0) := X"FF";
  CONSTANT CH1_B : STD_LOGIC_VECTOR(7 DOWNTO 0) := X"00";

  CONSTANT CH2_R : STD_LOGIC_VECTOR(7 DOWNTO 0) := X"00";
  CONSTANT CH2_G : STD_LOGIC_VECTOR(7 DOWNTO 0) := X"FF";
  CONSTANT CH2_B : STD_LOGIC_VECTOR(7 DOWNTO 0) := X"00";

  ----------------------------- STATES --------------------------------

  TYPE state_type IS (
    RESET_STATE,
    LONG_DELAY_STATE,
    RESET_AD7606_STATE,
    WAIT_FORCED_STATE,
    SET_STORE_FLAG_STATE,
    BEGIN_CONVERSION_STATE,
    ASSERT_CONVST_STATE,
    WAIT_BUSY_0_STATE,
    WAIT_BUSY_1_STATE,
    READ_CH1_LOW_STATE,
    WRITE_CH1_TRIGGER_STATE,
    WRITE_CH1_BRAM_STATE,
    READ_CH1_HIGH_STATE,
    RESET_SHORT_STATE,
    READ_CH2_LOW_STATE,
    WRITE_CH2_TRIGGER_STATE,
    WRITE_CH2_BRAM_STATE,
    READ_CH2_HIGH_STATE,
    WAIT_SAMPLE_INT_STATE,
    BRAM_FULL_STATE,
    CLEAR_STORE_FLAG_STATE
  );

  --- top level instantiations

  COMPONENT acquireToHDMI_fsm IS
  END COMPONENT;

  COMPONENT acquireToHDMI_datapath IS
    PORT (
      clk : IN STD_LOGIC;
      resetn : IN STD_LOGIC;
      cw : IN STD_LOGIC_VECTOR(CW_WIDTH - 1 DOWNTO 0);
      sw : OUT STD_LOGIC_VECTOR(DATAPATH_SW_WIDTH - 1 DOWNTO 0);
      an7606data : IN STD_LOGIC_VECTOR(15 DOWNTO 0);

      triggerVolt16bitSigned : IN SIGNED(15 DOWNTO 0);
      triggerTimePixel : IN STD_LOGIC_VECTOR(VIDEO_WIDTH_IN_BITS - 1 DOWNTO 0);
      ch1Data16bitSLV, ch2Data16bitSLV : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);

      tmdsDataP : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
      tmdsDataN : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
      tmdsClkP : OUT STD_LOGIC;
      tmdsClkN : OUT STD_LOGIC;
      hdmiOen : OUT STD_LOGIC
    );
  END COMPONENT;

  COMPONENT acquireToHDMI IS
  END COMPONENT;

  COMPONENT twosToPixel IS
    PORT (
      inputTwosComp : IN STD_LOGIC_VECTOR(16 DOWNTO 0),
      pixel : OUT STD_LOGIC_VECTOR(VIDEO_WIDTH_IN_BITS - 1 DOWNTO 0)
    );
  END COMPONENT;

  COMPONENT an7606 IS
    PORT (
      clk : IN STD_LOGIC;
      an7606data : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
      an7606convst, an7606cs, an7606rd, an7606reset : IN STD_LOGIC;
      an7606od : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      an7606busy : OUT STD_LOGIC);
  END COMPONENT;

  COMPONENT blk_mem_gen_0 IS
    PORT (
      clka : IN STD_LOGIC;
      ena : IN STD_LOGIC;
      wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      addra : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
      dina : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
      clkb : IN STD_LOGIC;
      enb : IN STD_LOGIC;
      addrb : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
      doutb : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
    );
  END COMPONENT;

END PACKAGE;