----------------------------------------------------------------------------------

----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.hdmi_package.all;


package acquireToHDMI_package is


-- Clock period definitions
CONSTANT clk_period : time := 20 ns;			-- 50Mhz crystal input (XTL_IN).

-- You need to complete this
type state_type is (RESET_STATE);


---------------------------- CONTROL WORD -----------------------------
CONSTANT CW_WIDTH : NATURAL := 22;
CONSTANT CONTROL_CW_WIDTH : NATURAL := xx;

CONSTANT CLEAR_STORE_FLAG_CW_BIT_INDEX : NATURAL := 21;
CONSTANT SET_STORE_FLAG_CW_BIT_INDEX : NATURAL := 20;
CONSTANT TRIG_CH2_WRITE_CW_BIT_INDEX : NATURAL := 19;
CONSTANT TRIG_CH1_WRITE_CW_BIT_INDEX : NATURAL := 18;
CONSTANT CONVERSION_PLUS_READOUT_CW_BIT_INDEX : NATURAL := 17;
CONSTANT SAMPLE_TIMER_ROLLOVER_CW_BIT_INDEX : NATURAL := 16;
CONSTANT DATA_STORAGE_CH2_WRITE_CW_BIT_INDEX : NATURAL := 15;
CONSTANT DATA_STORAGE_CH1_WRITE_CW_BIT_INDEX : NATURAL := 14;
CONSTANT CONVST_CW_BIT_INDEX : NATURAL := 13;
CONSTANT RD_CW_BIT_INDEX : NATURAL := 12;
CONSTANT CS_CW_BIT_INDEX : NATURAL := 11;
CONSTANT RESET_AD76076_CW_BIT_INDEX: NATURAL := 10;
CONSTANT DATA_STORAGE_COUNTER_CW_BIT1_INDEX : NATURAL := 9;
CONSTANT DATA_STORAGE_COUNTER_CW_BIT0_INDEX : NATURAL := 8;
CONSTANT SAMPLING_COUNTER_CW_BIT1_INDEX : NATURAL := 7;
CONSTANT SAMPLING_COUNTER_CW_BIT0_INDEX : NATURAL := 6;
CONSTANT SAMPLING_RATE_SELECT_CW_BIT1_INDEX : NATURAL := 5;
CONSTANT SAMPLING_RATE_SELECT_CW_BIT0_INDEX : NATURAL := 4;
CONSTANT LONG_DELAY_COUNTER_CW_BIT1_INDEX : NATURAL := 3;
CONSTANT LONG_DELAY_COUNTER_CW_BIT0_INDEX : NATURAL := 2;
CONSTANT SHORT_DELAY_COUNTER_CW_BIT1_INDEX : NATURAL := 1;
CONSTANT SHORT_DELAY_COUNTER_CW_BIT0_INDEX : NATURAL := 0;



---------------------------- STATUS WORD -----------------------------
CONSTANT SW_WIDTH : NATURAL := 12;
CONSTANT DATAPATH_SW_WIDTH : NATURAL := 6;

CONSTANT AD7606_BUSY_SW_INDEX :   NATURAL := 11;
CONSTANT STORE_TO_BRAM_SW_INDEX : NATURAL := 10;
CONSTANT CH2_TRIGGER_SW_INDEX :   NATURAL := 9;
CONSTANT CH1_TRIGGER_SW_INDEX :   NATURAL := 8;
CONSTANT LONG_DELAY_SW_INDEX :    NATURAL := 7;
CONSTANT SHORT_DELAY_SW_INDEX :   NATURAL := 6;
CONSTANT FULL_SW_INDEX :          NATURAL := 5;
CONSTANT SAMPLE_SW_INDEX :        NATURAL := 4;
CONSTANT TRIGGER_SW_INDEX :       NATURAL := 3;
CONSTANT STORE_SW_INDEX :         NATURAL := 2;
CONSTANT FORCED_SW_INDEX :        NATURAL := 1;
CONSTANT SINGLE_SW_INDEX :        NATURAL := 0;


------------------------- OTHER CONSTANTS ----------------------------

CONSTANT LONG_DELAY_50Mhz_CONST_WIDTH : NATURAL := 24;
CONSTANT LONG_DELAY_50Mhz_COUNTS : STD_LOGIC_VECTOR(LONG_DELAY_50Mhz_CONST_WIDTH - 1 downto 0) := x"00FFFF";

CONSTANT SHORT_DELAY_50Mhz_CONST_WIDTH : NATURAL := 8; 
CONSTANT SHORT_DELAY_50Mhz_COUNTS : STD_LOGIC_VECTOR(SHORT_DELAY_50Mhz_CONST_WIDTH - 1 downto 0) := x"10";

CONSTANT HIGHEST_RATE   : STD_LOGIC_VECTOR(31 downto 0) := STD_LOGIC_VECTOR(to_unsigned(300, 32));
CONSTANT HIGH_RATE      : STD_LOGIC_VECTOR(31 downto 0) := STD_LOGIC_VECTOR(to_unsigned(600, 32));
CONSTANT LOWEST_RATE    : STD_LOGIC_VECTOR(31 downto 0) := STD_LOGIC_VECTOR(to_unsigned(1200, 32));
CONSTANT LOW_RATE       : STD_LOGIC_VECTOR(31 downto 0) := STD_LOGIC_VECTOR(to_unsigned(2400, 32));

----------------------------- STATES --------------------------------

type state_type is (
  RESET_STATE,
  LONG_DELAY_STATE, 
  RESET_AD7606_STATE, 
  WAIT_FORCED_STATE,
  SET_STORE_FLAG_STATE,
  BEGIN_CONVERSION_STATE,
  ASSERT_CONVST_STATE,
  WAIT_BUSY_0_STATE, 
  WAIT_BUSY_1_STATE, 
  READ_CH1_LOW_STATE,
  WRITE_CH1_TRIGGER_STATE,
  WRITE_CH1_BRAM_STATE,
  READ_CH1_HIGH_STATE,        
  RESET_SHORT_STATE,
  READ_CH2_LOW_STATE,
  WRITE_CH2_TRIGGER_STATE,
  WRITE_CH2_BRAM_STATE,
  READ_CH2_HIGH_STATE,   
  WAIT_SAMPLE_INT_STATE, 
  BRAM_FULL_STATE,
  CLEAR_STORE_FLAG_STATE
  );

--- top level instantiations

component acquireToHDMI_fsm is
end component;

component acquireToHDMI_datapath is
end component;

component acquireToHDMI is
end component;	

component an7606 is
    PORT ( clk : in  STD_LOGIC;
           an7606data: out STD_LOGIC_VECTOR(15 downto 0);
           an7606convst, an7606cs, an7606rd, an7606reset: in STD_LOGIC;
           an7606od: in STD_LOGIC_VECTOR(2 downto 0);
           an7606busy : out STD_LOGIC);
END component;

component blk_mem_gen_0 is
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    clkb : IN STD_LOGIC;
    enb : IN STD_LOGIC;
    addrb : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    doutb : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
  );
END component;

end package;
